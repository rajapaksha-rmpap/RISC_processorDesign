library verilog;
use verilog.vl_types.all;
entity branch_tb is
end branch_tb;
