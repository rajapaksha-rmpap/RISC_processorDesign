library verilog;
use verilog.vl_types.all;
entity loadDataExt_tb is
end loadDataExt_tb;
