library verilog;
use verilog.vl_types.all;
entity pc_tb is
end pc_tb;
