library verilog;
use verilog.vl_types.all;
entity RISC_RV32I_cpu_tb is
end RISC_RV32I_cpu_tb;
