library verilog;
use verilog.vl_types.all;
entity test is
    port(
        \out\           : out    vl_logic
    );
end test;
